library verilog;
use verilog.vl_types.all;
entity frequencyDivider_vlg_vec_tst is
end frequencyDivider_vlg_vec_tst;
