library verilog;
use verilog.vl_types.all;
entity pulseGenerator_vlg_vec_tst is
end pulseGenerator_vlg_vec_tst;
