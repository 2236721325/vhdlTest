library verilog;
use verilog.vl_types.all;
entity RSTrigger_vlg_vec_tst is
end RSTrigger_vlg_vec_tst;
