library verilog;
use verilog.vl_types.all;
entity frequencyDivider_vlg_check_tst is
    port(
        clock_out       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end frequencyDivider_vlg_check_tst;
