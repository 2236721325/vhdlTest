library verilog;
use verilog.vl_types.all;
entity top_level_vlg_vec_tst is
end top_level_vlg_vec_tst;
