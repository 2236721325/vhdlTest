library verilog;
use verilog.vl_types.all;
entity digitalTube_vlg_vec_tst is
end digitalTube_vlg_vec_tst;
