library verilog;
use verilog.vl_types.all;
entity pulseGenerator_vlg_check_tst is
    port(
        fout            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end pulseGenerator_vlg_check_tst;
