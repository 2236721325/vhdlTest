library verilog;
use verilog.vl_types.all;
entity digitalCounter_vlg_vec_tst is
end digitalCounter_vlg_vec_tst;
