library verilog;
use verilog.vl_types.all;
entity fullAdderVector_vlg_vec_tst is
end fullAdderVector_vlg_vec_tst;
